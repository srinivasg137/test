module two_stage_sync(

);


endmodule